module vhumanise